/*
 * Copyright 2020 Google LLC
 * Copyright 2023 Frontgrade Gaisler
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *      http://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 */

// encoded as fmv instructions
`DEFINE_ZFA_INSTR(FLI_H,       I_FORMAT, ARITHMETIC, RV32ZFA);
`DEFINE_ZFA_INSTR(FLI_S,       I_FORMAT, ARITHMETIC, RV32ZFA);
`DEFINE_ZFA_INSTR(FLI_D,       I_FORMAT, ARITHMETIC, RV32ZFA);
`DEFINE_ZFA_INSTR(FLI_Q,       I_FORMAT, ARITHMETIC, RV32ZFA);
// encoded as fmin/fmax instructions
`DEFINE_ZFA_INSTR(FMINM_H,     R_FORMAT, ARITHMETIC, RV32ZFA);
`DEFINE_ZFA_INSTR(FMINM_S,     R_FORMAT, ARITHMETIC, RV32ZFA);
`DEFINE_ZFA_INSTR(FMINM_D,     R_FORMAT, ARITHMETIC, RV32ZFA);
`DEFINE_ZFA_INSTR(FMINM_Q,     R_FORMAT, ARITHMETIC, RV32ZFA);
`DEFINE_ZFA_INSTR(FMAXM_H,     R_FORMAT, ARITHMETIC, RV32ZFA);
`DEFINE_ZFA_INSTR(FMAXM_S,     R_FORMAT, ARITHMETIC, RV32ZFA);
`DEFINE_ZFA_INSTR(FMAXM_D,     R_FORMAT, ARITHMETIC, RV32ZFA);
`DEFINE_ZFA_INSTR(FMAXM_Q,     R_FORMAT, ARITHMETIC, RV32ZFA);
// encoded as fcvt
`DEFINE_ZFA_INSTR(FROUND_H,    I_FORMAT, ARITHMETIC, RV32ZFA);
`DEFINE_ZFA_INSTR(FROUNDNX_H,  I_FORMAT, ARITHMETIC, RV32ZFA);
`DEFINE_ZFA_INSTR(FROUND_S,    I_FORMAT, ARITHMETIC, RV32ZFA);
`DEFINE_ZFA_INSTR(FROUNDNX_S,  I_FORMAT, ARITHMETIC, RV32ZFA);
`DEFINE_ZFA_INSTR(FROUND_D,    I_FORMAT, ARITHMETIC, RV32ZFA);
`DEFINE_ZFA_INSTR(FROUNDNX_D,  I_FORMAT, ARITHMETIC, RV32ZFA);
`DEFINE_ZFA_INSTR(FROUND_Q,    I_FORMAT, ARITHMETIC, RV32ZFA);
`DEFINE_ZFA_INSTR(FROUNDNX_Q,  I_FORMAT, ARITHMETIC, RV32ZFA);
`DEFINE_ZFA_INSTR(FCVTMOD_W_D, I_FORMAT, ARITHMETIC, RV32ZFA);
`DEFINE_ZFA_INSTR(FMVH_X_D,    I_FORMAT, ARITHMETIC, RV32ZFA);
`DEFINE_ZFA_INSTR(FMVP_D_X,    R_FORMAT, ARITHMETIC, RV32ZFA);
// encoded as flt/fle...
`DEFINE_ZFA_INSTR(FLEQ_H,      R_FORMAT, COMPARE, RV32ZFA);
`DEFINE_ZFA_INSTR(FLTQ_H,      R_FORMAT, COMPARE, RV32ZFA);
`DEFINE_ZFA_INSTR(FLEQ_S,      R_FORMAT, COMPARE, RV32ZFA);
`DEFINE_ZFA_INSTR(FLTQ_S,      R_FORMAT, COMPARE, RV32ZFA);
`DEFINE_ZFA_INSTR(FLEQ_D,      R_FORMAT, COMPARE, RV32ZFA);
`DEFINE_ZFA_INSTR(FLTQ_D,      R_FORMAT, COMPARE, RV32ZFA);
`DEFINE_ZFA_INSTR(FLEQ_Q,      R_FORMAT, COMPARE, RV32ZFA);
`DEFINE_ZFA_INSTR(FLTQ_Q,      R_FORMAT, COMPARE, RV32ZFA);