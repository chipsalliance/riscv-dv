/*
 * Copyright 2020 Google LLC
 * Copyright 2023 Frontgrade Gaisler
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *      http://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 */

`DEFINE_FP_INSTR(FLH,       I_FORMAT,  LOAD,       RV32ZFH)
`DEFINE_FP_INSTR(FSH,       S_FORMAT,  STORE,      RV32ZFH)
`DEFINE_FP_INSTR(FMADD_H,   R4_FORMAT, ARITHMETIC, RV32ZFH)
`DEFINE_FP_INSTR(FMSUB_H,   R4_FORMAT, ARITHMETIC, RV32ZFH)
`DEFINE_FP_INSTR(FNMSUB_H,  R4_FORMAT, ARITHMETIC, RV32ZFH)
`DEFINE_FP_INSTR(FNMADD_H,  R4_FORMAT, ARITHMETIC, RV32ZFH)
`DEFINE_FP_INSTR(FADD_H,    R_FORMAT,  ARITHMETIC, RV32ZFH)
`DEFINE_FP_INSTR(FSUB_H,    R_FORMAT,  ARITHMETIC, RV32ZFH)
`DEFINE_FP_INSTR(FMUL_H,    R_FORMAT,  ARITHMETIC, RV32ZFH)
`DEFINE_FP_INSTR(FDIV_H,    R_FORMAT,  ARITHMETIC, RV32ZFH)
`DEFINE_FP_INSTR(FSQRT_H,   I_FORMAT,  ARITHMETIC, RV32ZFH)
`DEFINE_FP_INSTR(FSGNJ_H,   R_FORMAT,  ARITHMETIC, RV32ZFH)
`DEFINE_FP_INSTR(FSGNJN_H,  R_FORMAT,  ARITHMETIC, RV32ZFH)
`DEFINE_FP_INSTR(FSGNJX_H,  R_FORMAT,  ARITHMETIC, RV32ZFH)
`DEFINE_FP_INSTR(FMIN_H,    R_FORMAT,  ARITHMETIC, RV32ZFH)
`DEFINE_FP_INSTR(FMAX_H,    R_FORMAT,  ARITHMETIC, RV32ZFH)
`DEFINE_FP_INSTR(FCVT_S_H,  I_FORMAT,  ARITHMETIC, RV32ZFH)
`DEFINE_FP_INSTR(FCVT_H_S,  I_FORMAT,  ARITHMETIC, RV32ZFH)
`DEFINE_FP_INSTR(FCVT_D_H,  I_FORMAT,  ARITHMETIC, RV32ZFH)
`DEFINE_FP_INSTR(FCVT_H_D,  I_FORMAT,  ARITHMETIC, RV32ZFH)
`DEFINE_FP_INSTR(FCVT_Q_H,  I_FORMAT,  ARITHMETIC, RV32ZFH)
`DEFINE_FP_INSTR(FCVT_H_Q,  I_FORMAT,  ARITHMETIC, RV32ZFH)
`DEFINE_FP_INSTR(FEQ_H,     R_FORMAT,  COMPARE,    RV32ZFH)
`DEFINE_FP_INSTR(FLT_H,     R_FORMAT,  COMPARE,    RV32ZFH)
`DEFINE_FP_INSTR(FLE_H,     R_FORMAT,  COMPARE,    RV32ZFH)
`DEFINE_FP_INSTR(FCLASS_H,  R_FORMAT,  ARITHMETIC, RV32ZFH)
`DEFINE_FP_INSTR(FCVT_W_H,  I_FORMAT,  ARITHMETIC, RV32ZFH)
`DEFINE_FP_INSTR(FCVT_WU_H, I_FORMAT,  ARITHMETIC, RV32ZFH)
`DEFINE_FP_INSTR(FMV_X_H,   I_FORMAT,  ARITHMETIC, RV32ZFH)
`DEFINE_FP_INSTR(FCVT_H_W,  I_FORMAT,  ARITHMETIC, RV32ZFH)
`DEFINE_FP_INSTR(FCVT_H_WU, I_FORMAT,  ARITHMETIC, RV32ZFH)
`DEFINE_FP_INSTR(FMV_H_X,   I_FORMAT,  ARITHMETIC, RV32ZFH)
