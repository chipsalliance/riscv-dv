/*
 * Copyright 2020 Google LLC
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *      http://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 */

// Vector CSR access instruction
`DEFINE_INSTR(VSETVLI,    VSET_FORMAT, CSR, RV32V)
`DEFINE_INSTR(VSETVL,     VSET_FORMAT, CSR, RV32V)
// Vector integer arithmetic instruction
`DEFINE_VA_INSTR(VADD,     VA_FORMAT, ARITHMETIC, RV32V, {VV, VX, VI})
`DEFINE_VA_INSTR(VSUB,     VA_FORMAT, ARITHMETIC, RV32V, {VV, VX})
`DEFINE_VA_INSTR(VRSUB,    VA_FORMAT, ARITHMETIC, RV32V, {VX, VI})
`DEFINE_VA_INSTR(VWADDU,   VA_FORMAT, ARITHMETIC, RV32V, {VV, VX, WV, WX})
`DEFINE_VA_INSTR(VWSUBU,   VA_FORMAT, ARITHMETIC, RV32V, {VV, VX, WV, WX})
`DEFINE_VA_INSTR(VWADD,    VA_FORMAT, ARITHMETIC, RV32V, {VV, VX, WV, WX})
`DEFINE_VA_INSTR(VWSUB,    VA_FORMAT, ARITHMETIC, RV32V, {VV, VX, WV, WX})
`DEFINE_VA_INSTR(VADC,     VA_FORMAT, ARITHMETIC, RV32V, {VVM, VXM, VIM})
`DEFINE_VA_INSTR(VMADC,    VA_FORMAT, ARITHMETIC, RV32V, {VVM, VXM, VIM, VV, VX, VI})
`DEFINE_VA_INSTR(VSBC,     VA_FORMAT, ARITHMETIC, RV32V, {VVM, VXM})
`DEFINE_VA_INSTR(VMSBC,    VA_FORMAT, ARITHMETIC, RV32V, {VVM, VXM, VV, VX})
`DEFINE_VA_INSTR(VAND,     VA_FORMAT, ARITHMETIC, RV32V, {VV, VX, VI})
`DEFINE_VA_INSTR(VOR,      VA_FORMAT, ARITHMETIC, RV32V, {VV, VX, VI})
`DEFINE_VA_INSTR(VXOR,     VA_FORMAT, ARITHMETIC, RV32V, {VV, VX, VI})
`DEFINE_VA_INSTR(VSLL,     VA_FORMAT, SHIFT, RV32V, {VV, VX, VI})
`DEFINE_VA_INSTR(VSRL,     VA_FORMAT, SHIFT, RV32V, {VV, VX, VI})
`DEFINE_VA_INSTR(VSRA,     VA_FORMAT, SHIFT, RV32V, {VV, VX, VI})
`DEFINE_VA_INSTR(VNSRL,    VA_FORMAT, SHIFT, RV32V, {WV, WX, WI})
`DEFINE_VA_INSTR(VNSRA,    VA_FORMAT, SHIFT, RV32V, {WV, WX, WI})
`DEFINE_VA_INSTR(VMSEQ,    VA_FORMAT, COMPARE, RV32V, {VV, VX, VI})
`DEFINE_VA_INSTR(VMSNE,    VA_FORMAT, COMPARE, RV32V, {VV, VX, VI})
`DEFINE_VA_INSTR(VMSLTU,   VA_FORMAT, COMPARE, RV32V, {VV, VX})
`DEFINE_VA_INSTR(VMSLT,    VA_FORMAT, COMPARE, RV32V, {VV, VX})
`DEFINE_VA_INSTR(VMSLEU,   VA_FORMAT, COMPARE, RV32V, {VV, VX, VI})
`DEFINE_VA_INSTR(VMSLE,    VA_FORMAT, COMPARE, RV32V, {VV, VX, VI})
`DEFINE_VA_INSTR(VMSGTU,   VA_FORMAT, COMPARE, RV32V, {VX, VI})
`DEFINE_VA_INSTR(VMSGT,    VA_FORMAT, COMPARE, RV32V, {VX, VI})
`DEFINE_VA_INSTR(VMINU,    VA_FORMAT, ARITHMETIC, RV32V, {VV, VX})
`DEFINE_VA_INSTR(VMIN,     VA_FORMAT, ARITHMETIC, RV32V, {VV, VX})
`DEFINE_VA_INSTR(VMAXU,    VA_FORMAT, ARITHMETIC, RV32V, {VV, VX})
`DEFINE_VA_INSTR(VMAX,     VA_FORMAT, ARITHMETIC, RV32V, {VV, VX})
`DEFINE_VA_INSTR(VMUL,     VA_FORMAT, ARITHMETIC, RV32V, {VV, VX})
`DEFINE_VA_INSTR(VMULH,    VA_FORMAT, ARITHMETIC, RV32V, {VV, VX})
`DEFINE_VA_INSTR(VMULHU,   VA_FORMAT, ARITHMETIC, RV32V, {VV, VX})
`DEFINE_VA_INSTR(VMULHSU,  VA_FORMAT, ARITHMETIC, RV32V, {VV, VX})
`DEFINE_VA_INSTR(VDIVU,    VA_FORMAT, ARITHMETIC, RV32V, {VV, VX})
`DEFINE_VA_INSTR(VDIV,     VA_FORMAT, ARITHMETIC, RV32V, {VV, VX})
`DEFINE_VA_INSTR(VREMU,    VA_FORMAT, ARITHMETIC, RV32V, {VV, VX})
`DEFINE_VA_INSTR(VREM,     VA_FORMAT, ARITHMETIC, RV32V, {VV, VX})
`DEFINE_VA_INSTR(VWMUL,    VA_FORMAT, ARITHMETIC, RV32V, {VV, VX})
`DEFINE_VA_INSTR(VWMULU,   VA_FORMAT, ARITHMETIC, RV32V, {VV, VX})
`DEFINE_VA_INSTR(VWMULSU,  VA_FORMAT, ARITHMETIC, RV32V, {VV, VX})
`DEFINE_VA_INSTR(VMACC,    VA_FORMAT, ARITHMETIC, RV32V, {VV, VX})
`DEFINE_VA_INSTR(VNMSAC,   VA_FORMAT, ARITHMETIC, RV32V, {VV, VX})
`DEFINE_VA_INSTR(VMADD,    VA_FORMAT, ARITHMETIC, RV32V, {VV, VX})
`DEFINE_VA_INSTR(VNMSUB,   VA_FORMAT, ARITHMETIC, RV32V, {VV, VX})
`DEFINE_VA_INSTR(VWMACCU,  VA_FORMAT, ARITHMETIC, RV32V, {VV, VX})
`DEFINE_VA_INSTR(VWMACC,   VA_FORMAT, ARITHMETIC, RV32V, {VV, VX})
`DEFINE_VA_INSTR(VWMACCSU, VA_FORMAT, ARITHMETIC, RV32V, {VV, VX})
`DEFINE_VA_INSTR(VWMACCUS, VA_FORMAT, ARITHMETIC, RV32V, {VX})
/*
`DEFINE_VA_INSTR(VQMACCU,  VA_FORMAT, ARITHMETIC, RV32V, {VV, VX})
`DEFINE_VA_INSTR(VQMACC,   VA_FORMAT, ARITHMETIC, RV32V, {VV, VX})
`DEFINE_VA_INSTR(VQMACCSU, VA_FORMAT, ARITHMETIC, RV32V, {VV, VX})
`DEFINE_VA_INSTR(VQMACCUS, VA_FORMAT, ARITHMETIC, RV32V, {VX})
*/
`DEFINE_VA_INSTR(VMERGE,   VA_FORMAT, ARITHMETIC, RV32V, {VVM, VXM, VIM})
`DEFINE_VA_INSTR(VMV,      VA_FORMAT, ARITHMETIC, RV32V, {VV, VX, VI})
