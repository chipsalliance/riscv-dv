/*
 * Copyright 2020 Google LLC
 * Copyright 2023 Frontgrade Gaisler
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *      http://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 */

`DEFINE_ZFA_INSTR(FMVH_X_Q, I_FORMAT, ARITHMETIC, RV64ZFA);
`DEFINE_ZFA_INSTR(FMVP_Q_X, R_FORMAT, ARITHMETIC, RV64ZFA);
