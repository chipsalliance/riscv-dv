// Add your custom extensions, you can list all your local extended SV files here

`include "noelv_asm_program_gen.sv"