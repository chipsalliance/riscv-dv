
/*
 * Copyright 2020 Google LLC
 * Copyright 2023 Frontgrade Gaisler
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *      http://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 */

`DEFINE_FP_INSTR(FCVT_L_H,  I_FORMAT, ARITHMETIC, RV64ZFH)
`DEFINE_FP_INSTR(FCVT_LU_H, I_FORMAT, ARITHMETIC, RV64ZFH)
`DEFINE_FP_INSTR(FCVT_H_L,  I_FORMAT, ARITHMETIC, RV64ZFH)
`DEFINE_FP_INSTR(FCVT_H_LU, I_FORMAT, ARITHMETIC, RV64ZFH)
